module switch(
    //��λ�����Ѿ����ɣ��ڶ���ģ����ʵ��
    input clk,
    input [67:0] P_16,
    input [67:0] P_15,
    input [67:0] P_14,
    input [67:0] P_13,
    input [67:0] P_12,
    input [67:0] P_11,
    input [67:0] P_10,
    input [67:0] P_9,
    input [67:0] P_8,
    input [67:0] P_7,
    input [67:0] P_6,
    input [67:0] P_5,
    input [67:0] P_4,
    input [67:0] P_3,
    input [67:0] P_2,
    input [67:0] P_1,
    input [67:0] P_0,

    input c_16,
    input c_15,
    input c_14,
    input c_13,
    input c_12,
    input c_11,
    input c_10,
    input c_9,
    input c_8,
    input c_7,
    input c_6,
    input c_5,
    input c_4,
    input c_3,
    input c_2,
    input c_1,
    input c_0,

    output reg [16:0] c,
    output reg [16:0] In_wallace_0,
    output reg [16:0] In_wallace_1,
    output reg [16:0] In_wallace_2,
    output reg [16:0] In_wallace_3,
    output reg [16:0] In_wallace_4,
    output reg [16:0] In_wallace_5,
    output reg [16:0] In_wallace_6,
    output reg [16:0] In_wallace_7,
    output reg [16:0] In_wallace_8,
    output reg [16:0] In_wallace_9,
    output reg [16:0] In_wallace_10,
    output reg [16:0] In_wallace_11,
    output reg [16:0] In_wallace_12,
    output reg [16:0] In_wallace_13,
    output reg [16:0] In_wallace_14,
    output reg [16:0] In_wallace_15,
    output reg [16:0] In_wallace_16,
    output reg [16:0] In_wallace_17,
    output reg [16:0] In_wallace_18,
    output reg [16:0] In_wallace_19,
    output reg [16:0] In_wallace_20,
    output reg [16:0] In_wallace_21,
    output reg [16:0] In_wallace_22,
    output reg [16:0] In_wallace_23,
    output reg [16:0] In_wallace_24,
    output reg [16:0] In_wallace_25,
    output reg [16:0] In_wallace_26,
    output reg [16:0] In_wallace_27,
    output reg [16:0] In_wallace_28,
    output reg [16:0] In_wallace_29,
    output reg [16:0] In_wallace_30,
    output reg [16:0] In_wallace_31,
    output reg [16:0] In_wallace_32,
    output reg [16:0] In_wallace_33,
    output reg [16:0] In_wallace_34,
    output reg [16:0] In_wallace_35,
    output reg [16:0] In_wallace_36,
    output reg [16:0] In_wallace_37,
    output reg [16:0] In_wallace_38,
    output reg [16:0] In_wallace_39,
    output reg [16:0] In_wallace_40,
    output reg [16:0] In_wallace_41,
    output reg [16:0] In_wallace_42,
    output reg [16:0] In_wallace_43,
    output reg [16:0] In_wallace_44,
    output reg [16:0] In_wallace_45,
    output reg [16:0] In_wallace_46,
    output reg [16:0] In_wallace_47,
    output reg [16:0] In_wallace_48,
    output reg [16:0] In_wallace_49,
    output reg [16:0] In_wallace_50,
    output reg [16:0] In_wallace_51,
    output reg [16:0] In_wallace_52,
    output reg [16:0] In_wallace_53,
    output reg [16:0] In_wallace_54,
    output reg [16:0] In_wallace_55,
    output reg [16:0] In_wallace_56,
    output reg [16:0] In_wallace_57,
    output reg [16:0] In_wallace_58,
    output reg [16:0] In_wallace_59,
    output reg [16:0] In_wallace_60,
    output reg [16:0] In_wallace_61,
    output reg [16:0] In_wallace_62,
    output reg [16:0] In_wallace_63,
    output reg [16:0] In_wallace_64,
    output reg [16:0] In_wallace_65,
    output reg [16:0] In_wallace_66,
    output reg [16:0] In_wallace_67
);
always@(posedge clk)
begin
 c<={c_16,c_15,c_14,c_13,c_12,c_11,c_10,c_9,c_8,c_7,c_6,c_5,c_4,c_3,c_2,c_1,c_0};

 In_wallace_0<={P_16[0],P_15[0],P_14[0],P_13[0],P_12[0],P_11[0],P_10[0],P_9[0],P_8[0],P_7[0],P_6[0],P_5[0],P_4[0],P_3[0],P_2[0],P_1[0],P_0[0]};
 In_wallace_1<={P_16[1],P_15[1],P_14[1],P_13[1],P_12[1],P_11[1],P_10[1],P_9[1],P_8[1],P_7[1],P_6[1],P_5[1],P_4[1],P_3[1],P_2[1],P_1[1],P_0[1]};
 In_wallace_2<={P_16[2],P_15[2],P_14[2],P_13[2],P_12[2],P_11[2],P_10[2],P_9[2],P_8[2],P_7[2],P_6[2],P_5[2],P_4[2],P_3[2],P_2[2],P_1[2],P_0[2]};
 In_wallace_3<={P_16[3],P_15[3],P_14[3],P_13[3],P_12[3],P_11[3],P_10[3],P_9[3],P_8[3],P_7[3],P_6[3],P_5[3],P_4[3],P_3[3],P_2[3],P_1[3],P_0[3]};
 In_wallace_4<={P_16[4],P_15[4],P_14[4],P_13[4],P_12[4],P_11[4],P_10[4],P_9[4],P_8[4],P_7[4],P_6[4],P_5[4],P_4[4],P_3[4],P_2[4],P_1[4],P_0[4]};
 In_wallace_5<={P_16[5],P_15[5],P_14[5],P_13[5],P_12[5],P_11[5],P_10[5],P_9[5],P_8[5],P_7[5],P_6[5],P_5[5],P_4[5],P_3[5],P_2[5],P_1[5],P_0[5]};
 In_wallace_6<={P_16[6],P_15[6],P_14[6],P_13[6],P_12[6],P_11[6],P_10[6],P_9[6],P_8[6],P_7[6],P_6[6],P_5[6],P_4[6],P_3[6],P_2[6],P_1[6],P_0[6]};
 In_wallace_7<={P_16[7],P_15[7],P_14[7],P_13[7],P_12[7],P_11[7],P_10[7],P_9[7],P_8[7],P_7[7],P_6[7],P_5[7],P_4[7],P_3[7],P_2[7],P_1[7],P_0[7]};
 In_wallace_8<={P_16[8],P_15[8],P_14[8],P_13[8],P_12[8],P_11[8],P_10[8],P_9[8],P_8[8],P_7[8],P_6[8],P_5[8],P_4[8],P_3[8],P_2[8],P_1[8],P_0[8]};
 In_wallace_9<={P_16[9],P_15[9],P_14[9],P_13[9],P_12[9],P_11[9],P_10[9],P_9[9],P_8[9],P_7[9],P_6[9],P_5[9],P_4[9],P_3[9],P_2[9],P_1[9],P_0[9]};
 In_wallace_10<={P_16[10],P_15[10],P_14[10],P_13[10],P_12[10],P_11[10],P_10[10],P_9[10],P_8[10],P_7[10],P_6[10],P_5[10],P_4[10],P_3[10],P_2[10],P_1[10],P_0[10]};
 In_wallace_11<={P_16[11],P_15[11],P_14[11],P_13[11],P_12[11],P_11[11],P_10[11],P_9[11],P_8[11],P_7[11],P_6[11],P_5[11],P_4[11],P_3[11],P_2[11],P_1[11],P_0[11]};
 In_wallace_12<={P_16[12],P_15[12],P_14[12],P_13[12],P_12[12],P_11[12],P_10[12],P_9[12],P_8[12],P_7[12],P_6[12],P_5[12],P_4[12],P_3[12],P_2[12],P_1[12],P_0[12]};
 In_wallace_13<={P_16[13],P_15[13],P_14[13],P_13[13],P_12[13],P_11[13],P_10[13],P_9[13],P_8[13],P_7[13],P_6[13],P_5[13],P_4[13],P_3[13],P_2[13],P_1[13],P_0[13]};
 In_wallace_14<={P_16[14],P_15[14],P_14[14],P_13[14],P_12[14],P_11[14],P_10[14],P_9[14],P_8[14],P_7[14],P_6[14],P_5[14],P_4[14],P_3[14],P_2[14],P_1[14],P_0[14]};
 In_wallace_15<={P_16[15],P_15[15],P_14[15],P_13[15],P_12[15],P_11[15],P_10[15],P_9[15],P_8[15],P_7[15],P_6[15],P_5[15],P_4[15],P_3[15],P_2[15],P_1[15],P_0[15]};
     In_wallace_16<={P_16[16],P_15[16],P_14[16],P_13[16],P_12[16],P_11[16],P_10[16],P_9[16],P_8[16],P_7[16],P_6[16],P_5[16],P_4[16],P_3[16],P_2[16],P_1[16],P_0[16]};
     In_wallace_17<={P_16[17],P_15[17],P_14[17],P_13[17],P_12[17],P_11[17],P_10[17],P_9[17],P_8[17],P_7[17],P_6[17],P_5[17],P_4[17],P_3[17],P_2[17],P_1[17],P_0[17]};
     In_wallace_18<={P_16[18],P_15[18],P_14[18],P_13[18],P_12[18],P_11[18],P_10[18],P_9[18],P_8[18],P_7[18],P_6[18],P_5[18],P_4[18],P_3[18],P_2[18],P_1[18],P_0[18]};
     In_wallace_19<={P_16[19],P_15[19],P_14[19],P_13[19],P_12[19],P_11[19],P_10[19],P_9[19],P_8[19],P_7[19],P_6[19],P_5[19],P_4[19],P_3[19],P_2[19],P_1[19],P_0[19]};
     In_wallace_20<={P_16[20],P_15[20],P_14[20],P_13[20],P_12[20],P_11[20],P_10[20],P_9[20],P_8[20],P_7[20],P_6[20],P_5[20],P_4[20],P_3[20],P_2[20],P_1[20],P_0[20]};
     In_wallace_21<={P_16[21],P_15[21],P_14[21],P_13[21],P_12[21],P_11[21],P_10[21],P_9[21],P_8[21],P_7[21],P_6[21],P_5[21],P_4[21],P_3[21],P_2[21],P_1[21],P_0[21]};
     In_wallace_22<={P_16[22],P_15[22],P_14[22],P_13[22],P_12[22],P_11[22],P_10[22],P_9[22],P_8[22],P_7[22],P_6[22],P_5[22],P_4[22],P_3[22],P_2[22],P_1[22],P_0[22]};
     In_wallace_23<={P_16[23],P_15[23],P_14[23],P_13[23],P_12[23],P_11[23],P_10[23],P_9[23],P_8[23],P_7[23],P_6[23],P_5[23],P_4[23],P_3[23],P_2[23],P_1[23],P_0[23]};
     In_wallace_24<={P_16[24],P_15[24],P_14[24],P_13[24],P_12[24],P_11[24],P_10[24],P_9[24],P_8[24],P_7[24],P_6[24],P_5[24],P_4[24],P_3[24],P_2[24],P_1[24],P_0[24]};
     In_wallace_25<={P_16[25],P_15[25],P_14[25],P_13[25],P_12[25],P_11[25],P_10[25],P_9[25],P_8[25],P_7[25],P_6[25],P_5[25],P_4[25],P_3[25],P_2[25],P_1[25],P_0[25]};
     In_wallace_26<={P_16[26],P_15[26],P_14[26],P_13[26],P_12[26],P_11[26],P_10[26],P_9[26],P_8[26],P_7[26],P_6[26],P_5[26],P_4[26],P_3[26],P_2[26],P_1[26],P_0[26]};
     In_wallace_27<={P_16[27],P_15[27],P_14[27],P_13[27],P_12[27],P_11[27],P_10[27],P_9[27],P_8[27],P_7[27],P_6[27],P_5[27],P_4[27],P_3[27],P_2[27],P_1[27],P_0[27]};
     In_wallace_28<={P_16[28],P_15[28],P_14[28],P_13[28],P_12[28],P_11[28],P_10[28],P_9[28],P_8[28],P_7[28],P_6[28],P_5[28],P_4[28],P_3[28],P_2[28],P_1[28],P_0[28]};
     In_wallace_29<={P_16[29],P_15[29],P_14[29],P_13[29],P_12[29],P_11[29],P_10[29],P_9[29],P_8[29],P_7[29],P_6[29],P_5[29],P_4[29],P_3[29],P_2[29],P_1[29],P_0[29]};
     In_wallace_30<={P_16[30],P_15[30],P_14[30],P_13[30],P_12[30],P_11[30],P_10[30],P_9[30],P_8[30],P_7[30],P_6[30],P_5[30],P_4[30],P_3[30],P_2[30],P_1[30],P_0[30]};
     In_wallace_31<={P_16[31],P_15[31],P_14[31],P_13[31],P_12[31],P_11[31],P_10[31],P_9[31],P_8[31],P_7[31],P_6[31],P_5[31],P_4[31],P_3[31],P_2[31],P_1[31],P_0[31]};
     In_wallace_32<={P_16[32],P_15[32],P_14[32],P_13[32],P_12[32],P_11[32],P_10[32],P_9[32],P_8[32],P_7[32],P_6[32],P_5[32],P_4[32],P_3[32],P_2[32],P_1[32],P_0[32]};
     In_wallace_33<={P_16[33],P_15[33],P_14[33],P_13[33],P_12[33],P_11[33],P_10[33],P_9[33],P_8[33],P_7[33],P_6[33],P_5[33],P_4[33],P_3[33],P_2[33],P_1[33],P_0[33]};
     In_wallace_34<={P_16[34],P_15[34],P_14[34],P_13[34],P_12[34],P_11[34],P_10[34],P_9[34],P_8[34],P_7[34],P_6[34],P_5[34],P_4[34],P_3[34],P_2[34],P_1[34],P_0[34]};
     In_wallace_35<={P_16[35],P_15[35],P_14[35],P_13[35],P_12[35],P_11[35],P_10[35],P_9[35],P_8[35],P_7[35],P_6[35],P_5[35],P_4[35],P_3[35],P_2[35],P_1[35],P_0[35]};
     In_wallace_36<={P_16[36],P_15[36],P_14[36],P_13[36],P_12[36],P_11[36],P_10[36],P_9[36],P_8[36],P_7[36],P_6[36],P_5[36],P_4[36],P_3[36],P_2[36],P_1[36],P_0[36]};
     In_wallace_37<={P_16[37],P_15[37],P_14[37],P_13[37],P_12[37],P_11[37],P_10[37],P_9[37],P_8[37],P_7[37],P_6[37],P_5[37],P_4[37],P_3[37],P_2[37],P_1[37],P_0[37]};
     In_wallace_38<={P_16[38],P_15[38],P_14[38],P_13[38],P_12[38],P_11[38],P_10[38],P_9[38],P_8[38],P_7[38],P_6[38],P_5[38],P_4[38],P_3[38],P_2[38],P_1[38],P_0[38]};
     In_wallace_39<={P_16[39],P_15[39],P_14[39],P_13[39],P_12[39],P_11[39],P_10[39],P_9[39],P_8[39],P_7[39],P_6[39],P_5[39],P_4[39],P_3[39],P_2[39],P_1[39],P_0[39]};
     In_wallace_40<={P_16[40],P_15[40],P_14[40],P_13[40],P_12[40],P_11[40],P_10[40],P_9[40],P_8[40],P_7[40],P_6[40],P_5[40],P_4[40],P_3[40],P_2[40],P_1[40],P_0[40]};
     In_wallace_41<={P_16[41],P_15[41],P_14[41],P_13[41],P_12[41],P_11[41],P_10[41],P_9[41],P_8[41],P_7[41],P_6[41],P_5[41],P_4[41],P_3[41],P_2[41],P_1[41],P_0[41]};
     In_wallace_42<={P_16[42],P_15[42],P_14[42],P_13[42],P_12[42],P_11[42],P_10[42],P_9[42],P_8[42],P_7[42],P_6[42],P_5[42],P_4[42],P_3[42],P_2[42],P_1[42],P_0[42]};
     In_wallace_43<={P_16[43],P_15[43],P_14[43],P_13[43],P_12[43],P_11[43],P_10[43],P_9[43],P_8[43],P_7[43],P_6[43],P_5[43],P_4[43],P_3[43],P_2[43],P_1[43],P_0[43]};
     In_wallace_44<={P_16[44],P_15[44],P_14[44],P_13[44],P_12[44],P_11[44],P_10[44],P_9[44],P_8[44],P_7[44],P_6[44],P_5[44],P_4[44],P_3[44],P_2[44],P_1[44],P_0[44]};
     In_wallace_45<={P_16[45],P_15[45],P_14[45],P_13[45],P_12[45],P_11[45],P_10[45],P_9[45],P_8[45],P_7[45],P_6[45],P_5[45],P_4[45],P_3[45],P_2[45],P_1[45],P_0[45]};
     In_wallace_46<={P_16[46],P_15[46],P_14[46],P_13[46],P_12[46],P_11[46],P_10[46],P_9[46],P_8[46],P_7[46],P_6[46],P_5[46],P_4[46],P_3[46],P_2[46],P_1[46],P_0[46]};
     In_wallace_47<={P_16[47],P_15[47],P_14[47],P_13[47],P_12[47],P_11[47],P_10[47],P_9[47],P_8[47],P_7[47],P_6[47],P_5[47],P_4[47],P_3[47],P_2[47],P_1[47],P_0[47]};
     In_wallace_48<={P_16[48],P_15[48],P_14[48],P_13[48],P_12[48],P_11[48],P_10[48],P_9[48],P_8[48],P_7[48],P_6[48],P_5[48],P_4[48],P_3[48],P_2[48],P_1[48],P_0[48]};
     In_wallace_49<={P_16[49],P_15[49],P_14[49],P_13[49],P_12[49],P_11[49],P_10[49],P_9[49],P_8[49],P_7[49],P_6[49],P_5[49],P_4[49],P_3[49],P_2[49],P_1[49],P_0[49]};
     In_wallace_50<={P_16[50],P_15[50],P_14[50],P_13[50],P_12[50],P_11[50],P_10[50],P_9[50],P_8[50],P_7[50],P_6[50],P_5[50],P_4[50],P_3[50],P_2[50],P_1[50],P_0[50]};
     In_wallace_51<={P_16[51],P_15[51],P_14[51],P_13[51],P_12[51],P_11[51],P_10[51],P_9[51],P_8[51],P_7[51],P_6[51],P_5[51],P_4[51],P_3[51],P_2[51],P_1[51],P_0[51]};
     In_wallace_52<={P_16[52],P_15[52],P_14[52],P_13[52],P_12[52],P_11[52],P_10[52],P_9[52],P_8[52],P_7[52],P_6[52],P_5[52],P_4[52],P_3[52],P_2[52],P_1[52],P_0[52]};
     In_wallace_53<={P_16[53],P_15[53],P_14[53],P_13[53],P_12[53],P_11[53],P_10[53],P_9[53],P_8[53],P_7[53],P_6[53],P_5[53],P_4[53],P_3[53],P_2[53],P_1[53],P_0[53]};
     In_wallace_54<={P_16[54],P_15[54],P_14[54],P_13[54],P_12[54],P_11[54],P_10[54],P_9[54],P_8[54],P_7[54],P_6[54],P_5[54],P_4[54],P_3[54],P_2[54],P_1[54],P_0[54]};
     In_wallace_55<={P_16[55],P_15[55],P_14[55],P_13[55],P_12[55],P_11[55],P_10[55],P_9[55],P_8[55],P_7[55],P_6[55],P_5[55],P_4[55],P_3[55],P_2[55],P_1[55],P_0[55]};
     In_wallace_56<={P_16[56],P_15[56],P_14[56],P_13[56],P_12[56],P_11[56],P_10[56],P_9[56],P_8[56],P_7[56],P_6[56],P_5[56],P_4[56],P_3[56],P_2[56],P_1[56],P_0[56]};
     In_wallace_57<={P_16[57],P_15[57],P_14[57],P_13[57],P_12[57],P_11[57],P_10[57],P_9[57],P_8[57],P_7[57],P_6[57],P_5[57],P_4[57],P_3[57],P_2[57],P_1[57],P_0[57]};
     In_wallace_58<={P_16[58],P_15[58],P_14[58],P_13[58],P_12[58],P_11[58],P_10[58],P_9[58],P_8[58],P_7[58],P_6[58],P_5[58],P_4[58],P_3[58],P_2[58],P_1[58],P_0[58]};
     In_wallace_59<={P_16[59],P_15[59],P_14[59],P_13[59],P_12[59],P_11[59],P_10[59],P_9[59],P_8[59],P_7[59],P_6[59],P_5[59],P_4[59],P_3[59],P_2[59],P_1[59],P_0[59]};
     In_wallace_60<={P_16[60],P_15[60],P_14[60],P_13[60],P_12[60],P_11[60],P_10[60],P_9[60],P_8[60],P_7[60],P_6[60],P_5[60],P_4[60],P_3[60],P_2[60],P_1[60],P_0[60]};
     In_wallace_61<={P_16[61],P_15[61],P_14[61],P_13[61],P_12[61],P_11[61],P_10[61],P_9[61],P_8[61],P_7[61],P_6[61],P_5[61],P_4[61],P_3[61],P_2[61],P_1[61],P_0[61]};
     In_wallace_62<={P_16[62],P_15[62],P_14[62],P_13[62],P_12[62],P_11[62],P_10[62],P_9[62],P_8[62],P_7[62],P_6[62],P_5[62],P_4[62],P_3[62],P_2[62],P_1[62],P_0[62]};
     In_wallace_63<={P_16[63],P_15[63],P_14[63],P_13[63],P_12[63],P_11[63],P_10[63],P_9[63],P_8[63],P_7[63],P_6[63],P_5[63],P_4[63],P_3[63],P_2[63],P_1[63],P_0[63]};
     In_wallace_64<={P_16[64],P_15[64],P_14[64],P_13[64],P_12[64],P_11[64],P_10[64],P_9[64],P_8[64],P_7[64],P_6[64],P_5[64],P_4[64],P_3[64],P_2[64],P_1[64],P_0[64]};
     In_wallace_65<={P_16[65],P_15[65],P_14[65],P_13[65],P_12[65],P_11[65],P_10[65],P_9[65],P_8[65],P_7[65],P_6[65],P_5[65],P_4[65],P_3[65],P_2[65],P_1[65],P_0[65]};
     In_wallace_66<={P_16[66],P_15[66],P_14[66],P_13[66],P_12[66],P_11[66],P_10[66],P_9[66],P_8[66],P_7[66],P_6[66],P_5[66],P_4[66],P_3[66],P_2[66],P_1[66],P_0[66]};
     In_wallace_67<={P_16[67],P_15[67],P_14[67],P_13[67],P_12[67],P_11[67],P_10[67],P_9[67],P_8[67],P_7[67],P_6[67],P_5[67],P_4[67],P_3[67],P_2[67],P_1[67],P_0[67]};


end
    endmodule